// sdram.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module sdram (
		input  wire        clk_clk,             //   clk.clk
		input  wire        reset_reset_n,       // reset.reset_n
		input  wire [24:0] sdram_address,       // sdram.address
		input  wire [1:0]  sdram_byteenable_n,  //      .byteenable_n
		input  wire        sdram_chipselect,    //      .chipselect
		input  wire [15:0] sdram_writedata,     //      .writedata
		input  wire        sdram_read_n,        //      .read_n
		input  wire        sdram_write_n,       //      .write_n
		output wire [15:0] sdram_readdata,      //      .readdata
		output wire        sdram_readdatavalid, //      .readdatavalid
		output wire        sdram_waitrequest,   //      .waitrequest
		output wire [12:0] wire_addr,           //  wire.addr
		output wire [1:0]  wire_ba,             //      .ba
		output wire        wire_cas_n,          //      .cas_n
		output wire        wire_cke,            //      .cke
		output wire        wire_cs_n,           //      .cs_n
		inout  wire [15:0] wire_dq,             //      .dq
		output wire [1:0]  wire_dqm,            //      .dqm
		output wire        wire_ras_n,          //      .ras_n
		output wire        wire_we_n            //      .we_n
	);

	wire    sys_sdram_pll_0_sys_clk_clk;    // sys_sdram_pll_0:sys_clk_clk -> [new_sdram_controller_0:clk, rst_controller:clk]
	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> new_sdram_controller_0:reset_n

	sdram_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),     //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset), // reset.reset_n
		.az_addr        (sdram_address),                   //    s1.address
		.az_be_n        (sdram_byteenable_n),              //      .byteenable_n
		.az_cs          (sdram_chipselect),                //      .chipselect
		.az_data        (sdram_writedata),                 //      .writedata
		.az_rd_n        (sdram_read_n),                    //      .read_n
		.az_wr_n        (sdram_write_n),                   //      .write_n
		.za_data        (sdram_readdata),                  //      .readdata
		.za_valid       (sdram_readdatavalid),             //      .readdatavalid
		.za_waitrequest (sdram_waitrequest),               //      .waitrequest
		.zs_addr        (wire_addr),                       //  wire.export
		.zs_ba          (wire_ba),                         //      .export
		.zs_cas_n       (wire_cas_n),                      //      .export
		.zs_cke         (wire_cke),                        //      .export
		.zs_cs_n        (wire_cs_n),                       //      .export
		.zs_dq          (wire_dq),                         //      .export
		.zs_dqm         (wire_dqm),                        //      .export
		.zs_ras_n       (wire_ras_n),                      //      .export
		.zs_we_n        (wire_we_n)                        //      .export
	);

	sdram_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                     //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),              //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk), //      sys_clk.clk
		.sdram_clk_clk      (),                            //    sdram_clk.clk
		.reset_source_reset ()                             // reset_source.reset
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
